`ifndef _constants_vh_
`define _constants_vh_

`define nBits 264
`define nSBox 33

`define INIT_SBOX_LAYER\
		sBoxLayer[0] = 8'hee;	sBoxLayer[1] = 8'hed;	sBoxLayer[2] = 8'heb;	sBoxLayer[3] = 8'he0;	sBoxLayer[4] = 8'he2;	sBoxLayer[5] = 8'he1;	sBoxLayer[6] = 8'he4;	sBoxLayer[7] = 8'hef;	sBoxLayer[8] = 8'he7;	sBoxLayer[9] = 8'hea;	sBoxLayer[10] = 8'he8;	sBoxLayer[11] = 8'he5;	sBoxLayer[12] = 8'he9;	sBoxLayer[13] = 8'hec;	sBoxLayer[14] = 8'he3;	sBoxLayer[15] = 8'he6;\
		sBoxLayer[16] = 8'hde;	sBoxLayer[17] = 8'hdd;	sBoxLayer[18] = 8'hdb;	sBoxLayer[19] = 8'hd0;	sBoxLayer[20] = 8'hd2;	sBoxLayer[21] = 8'hd1;	sBoxLayer[22] = 8'hd4;	sBoxLayer[23] = 8'hdf;	sBoxLayer[24] = 8'hd7;	sBoxLayer[25] = 8'hda;	sBoxLayer[26] = 8'hd8;	sBoxLayer[27] = 8'hd5;	sBoxLayer[28] = 8'hd9;	sBoxLayer[29] = 8'hdc;	sBoxLayer[30] = 8'hd3;	sBoxLayer[31] = 8'hd6;\
		sBoxLayer[32] = 8'hbe;	sBoxLayer[33] = 8'hbd;	sBoxLayer[34] = 8'hbb;	sBoxLayer[35] = 8'hb0;	sBoxLayer[36] = 8'hb2;	sBoxLayer[37] = 8'hb1;	sBoxLayer[38] = 8'hb4;	sBoxLayer[39] = 8'hbf;	sBoxLayer[40] = 8'hb7;	sBoxLayer[41] = 8'hba;	sBoxLayer[42] = 8'hb8;	sBoxLayer[43] = 8'hb5;	sBoxLayer[44] = 8'hb9;	sBoxLayer[45] = 8'hbc;	sBoxLayer[46] = 8'hb3;	sBoxLayer[47] = 8'hb6;\
		sBoxLayer[48] = 8'h0e;	sBoxLayer[49] = 8'h0d;	sBoxLayer[50] = 8'h0b;	sBoxLayer[51] = 8'h00;	sBoxLayer[52] = 8'h02;	sBoxLayer[53] = 8'h01;	sBoxLayer[54] = 8'h04;	sBoxLayer[55] = 8'h0f;	sBoxLayer[56] = 8'h07;	sBoxLayer[57] = 8'h0a;	sBoxLayer[58] = 8'h08;	sBoxLayer[59] = 8'h05;	sBoxLayer[60] = 8'h09;	sBoxLayer[61] = 8'h0c;	sBoxLayer[62] = 8'h03;	sBoxLayer[63] = 8'h06;\
		sBoxLayer[64] = 8'h2e;	sBoxLayer[65] = 8'h2d;	sBoxLayer[66] = 8'h2b;	sBoxLayer[67] = 8'h20;	sBoxLayer[68] = 8'h22;	sBoxLayer[69] = 8'h21;	sBoxLayer[70] = 8'h24;	sBoxLayer[71] = 8'h2f;	sBoxLayer[72] = 8'h27;	sBoxLayer[73] = 8'h2a;	sBoxLayer[74] = 8'h28;	sBoxLayer[75] = 8'h25;	sBoxLayer[76] = 8'h29;	sBoxLayer[77] = 8'h2c;	sBoxLayer[78] = 8'h23;	sBoxLayer[79] = 8'h26;\
		sBoxLayer[80] = 8'h1e;	sBoxLayer[81] = 8'h1d;	sBoxLayer[82] = 8'h1b;	sBoxLayer[83] = 8'h10;	sBoxLayer[84] = 8'h12;	sBoxLayer[85] = 8'h11;	sBoxLayer[86] = 8'h14;	sBoxLayer[87] = 8'h1f;	sBoxLayer[88] = 8'h17;	sBoxLayer[89] = 8'h1a;	sBoxLayer[90] = 8'h18;	sBoxLayer[91] = 8'h15;	sBoxLayer[92] = 8'h19;	sBoxLayer[93] = 8'h1c;	sBoxLayer[94] = 8'h13;	sBoxLayer[95] = 8'h16;\
		sBoxLayer[96] = 8'h4e;	sBoxLayer[97] = 8'h4d;	sBoxLayer[98] = 8'h4b;	sBoxLayer[99] = 8'h40;	sBoxLayer[100] = 8'h42;	sBoxLayer[101] = 8'h41;	sBoxLayer[102] = 8'h44;	sBoxLayer[103] = 8'h4f;	sBoxLayer[104] = 8'h47;	sBoxLayer[105] = 8'h4a;	sBoxLayer[106] = 8'h48;	sBoxLayer[107] = 8'h45;	sBoxLayer[108] = 8'h49;	sBoxLayer[109] = 8'h4c;	sBoxLayer[110] = 8'h43;	sBoxLayer[111] = 8'h46;\
		sBoxLayer[112] = 8'hfe;	sBoxLayer[113] = 8'hfd;	sBoxLayer[114] = 8'hfb;	sBoxLayer[115] = 8'hf0;	sBoxLayer[116] = 8'hf2;	sBoxLayer[117] = 8'hf1;	sBoxLayer[118] = 8'hf4;	sBoxLayer[119] = 8'hff;	sBoxLayer[120] = 8'hf7;	sBoxLayer[121] = 8'hfa;	sBoxLayer[122] = 8'hf8;	sBoxLayer[123] = 8'hf5;	sBoxLayer[124] = 8'hf9;	sBoxLayer[125] = 8'hfc;	sBoxLayer[126] = 8'hf3;	sBoxLayer[127] = 8'hf6;\
		sBoxLayer[128] = 8'h7e;	sBoxLayer[129] = 8'h7d;	sBoxLayer[130] = 8'h7b;	sBoxLayer[131] = 8'h70;	sBoxLayer[132] = 8'h72;	sBoxLayer[133] = 8'h71;	sBoxLayer[134] = 8'h74;	sBoxLayer[135] = 8'h7f;	sBoxLayer[136] = 8'h77;	sBoxLayer[137] = 8'h7a;	sBoxLayer[138] = 8'h78;	sBoxLayer[139] = 8'h75;	sBoxLayer[140] = 8'h79;	sBoxLayer[141] = 8'h7c;	sBoxLayer[142] = 8'h73;	sBoxLayer[143] = 8'h76;\
		sBoxLayer[144] = 8'hae;	sBoxLayer[145] = 8'had;	sBoxLayer[146] = 8'hab;	sBoxLayer[147] = 8'ha0;	sBoxLayer[148] = 8'ha2;	sBoxLayer[149] = 8'ha1;	sBoxLayer[150] = 8'ha4;	sBoxLayer[151] = 8'haf;	sBoxLayer[152] = 8'ha7;	sBoxLayer[153] = 8'haa;	sBoxLayer[154] = 8'ha8;	sBoxLayer[155] = 8'ha5;	sBoxLayer[156] = 8'ha9;	sBoxLayer[157] = 8'hac;	sBoxLayer[158] = 8'ha3;	sBoxLayer[159] = 8'ha6;\
		sBoxLayer[160] = 8'h8e;	sBoxLayer[161] = 8'h8d;	sBoxLayer[162] = 8'h8b;	sBoxLayer[163] = 8'h80;	sBoxLayer[164] = 8'h82;	sBoxLayer[165] = 8'h81;	sBoxLayer[166] = 8'h84;	sBoxLayer[167] = 8'h8f;	sBoxLayer[168] = 8'h87;	sBoxLayer[169] = 8'h8a;	sBoxLayer[170] = 8'h88;	sBoxLayer[171] = 8'h85;	sBoxLayer[172] = 8'h89;	sBoxLayer[173] = 8'h8c;	sBoxLayer[174] = 8'h83;	sBoxLayer[175] = 8'h86;\
		sBoxLayer[176] = 8'h5e;	sBoxLayer[177] = 8'h5d;	sBoxLayer[178] = 8'h5b;	sBoxLayer[179] = 8'h50;	sBoxLayer[180] = 8'h52;	sBoxLayer[181] = 8'h51;	sBoxLayer[182] = 8'h54;	sBoxLayer[183] = 8'h5f;	sBoxLayer[184] = 8'h57;	sBoxLayer[185] = 8'h5a;	sBoxLayer[186] = 8'h58;	sBoxLayer[187] = 8'h55;	sBoxLayer[188] = 8'h59;	sBoxLayer[189] = 8'h5c;	sBoxLayer[190] = 8'h53;	sBoxLayer[191] = 8'h56;\
		sBoxLayer[192] = 8'h9e;	sBoxLayer[193] = 8'h9d;	sBoxLayer[194] = 8'h9b;	sBoxLayer[195] = 8'h90;	sBoxLayer[196] = 8'h92;	sBoxLayer[197] = 8'h91;	sBoxLayer[198] = 8'h94;	sBoxLayer[199] = 8'h9f;	sBoxLayer[200] = 8'h97;	sBoxLayer[201] = 8'h9a;	sBoxLayer[202] = 8'h98;	sBoxLayer[203] = 8'h95;	sBoxLayer[204] = 8'h99;	sBoxLayer[205] = 8'h9c;	sBoxLayer[206] = 8'h93;	sBoxLayer[207] = 8'h96;\
		sBoxLayer[208] = 8'hce;	sBoxLayer[209] = 8'hcd;	sBoxLayer[210] = 8'hcb;	sBoxLayer[211] = 8'hc0;	sBoxLayer[212] = 8'hc2;	sBoxLayer[213] = 8'hc1;	sBoxLayer[214] = 8'hc4;	sBoxLayer[215] = 8'hcf;	sBoxLayer[216] = 8'hc7;	sBoxLayer[217] = 8'hca;	sBoxLayer[218] = 8'hc8;	sBoxLayer[219] = 8'hc5;	sBoxLayer[220] = 8'hc9;	sBoxLayer[221] = 8'hcc;	sBoxLayer[222] = 8'hc3;	sBoxLayer[223] = 8'hc6;\
		sBoxLayer[224] = 8'h3e;	sBoxLayer[225] = 8'h3d;	sBoxLayer[226] = 8'h3b;	sBoxLayer[227] = 8'h30;	sBoxLayer[228] = 8'h32;	sBoxLayer[229] = 8'h31;	sBoxLayer[230] = 8'h34;	sBoxLayer[231] = 8'h3f;	sBoxLayer[232] = 8'h37;	sBoxLayer[233] = 8'h3a;	sBoxLayer[234] = 8'h38;	sBoxLayer[235] = 8'h35;	sBoxLayer[236] = 8'h39;	sBoxLayer[237] = 8'h3c;	sBoxLayer[238] = 8'h33;	sBoxLayer[239] = 8'h36;\
		sBoxLayer[240] = 8'h6e;	sBoxLayer[241] = 8'h6d;	sBoxLayer[242] = 8'h6b;	sBoxLayer[243] = 8'h60;	sBoxLayer[244] = 8'h62;	sBoxLayer[245] = 8'h61;	sBoxLayer[246] = 8'h64;	sBoxLayer[247] = 8'h6f;	sBoxLayer[248] = 8'h67;	sBoxLayer[249] = 8'h6a;	sBoxLayer[250] = 8'h68;	sBoxLayer[251] = 8'h65;	sBoxLayer[252] = 8'h69;	sBoxLayer[253] = 8'h6c;	sBoxLayer[254] = 8'h63;	sBoxLayer[255] = 8'h66;
`endif
