`ifndef _constants_vh_
`define _constants_vh_

`define nBits 264
`define nSBox 33

`endif
