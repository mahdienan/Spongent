`ifndef _constants_vh_
`define _constants_vh_

`define nBits 264				// = (capacity + rate) = (176 + 88)
`define nSBox 33				// = (nBits / 8) = (264 / 8)
`define rate 88
`define R_SizeInBytes 11 	// = (rate / 8) = (88 / 8)
`define nRounds 135

`define INIT_SBOX_LAYER\
sBoxLayer[0+:8] = 8'hee;\
sBoxLayer[8+:8] = 8'hed;\
sBoxLayer[16+:8] = 8'heb;\
sBoxLayer[24+:8] = 8'he0;\
sBoxLayer[32+:8] = 8'he2;\
sBoxLayer[40+:8] = 8'he1;\
sBoxLayer[48+:8] = 8'he4;\
sBoxLayer[56+:8] = 8'hef;\
sBoxLayer[64+:8] = 8'he7;\
sBoxLayer[72+:8] = 8'hea;\
sBoxLayer[80+:8] = 8'he8;\
sBoxLayer[88+:8] = 8'he5;\
sBoxLayer[96+:8] = 8'he9;\
sBoxLayer[104+:8] = 8'hec;\
sBoxLayer[112+:8] = 8'he3;\
sBoxLayer[120+:8] = 8'he6;\
sBoxLayer[128+:8] = 8'hde;\
sBoxLayer[136+:8] = 8'hdd;\
sBoxLayer[144+:8] = 8'hdb;\
sBoxLayer[152+:8] = 8'hd0;\
sBoxLayer[160+:8] = 8'hd2;\
sBoxLayer[168+:8] = 8'hd1;\
sBoxLayer[176+:8] = 8'hd4;\
sBoxLayer[184+:8] = 8'hdf;\
sBoxLayer[192+:8] = 8'hd7;\
sBoxLayer[200+:8] = 8'hda;\
sBoxLayer[208+:8] = 8'hd8;\
sBoxLayer[216+:8] = 8'hd5;\
sBoxLayer[224+:8] = 8'hd9;\
sBoxLayer[232+:8] = 8'hdc;\
sBoxLayer[240+:8] = 8'hd3;\
sBoxLayer[248+:8] = 8'hd6;\
sBoxLayer[256+:8] = 8'hbe;\
sBoxLayer[264+:8] = 8'hbd;\
sBoxLayer[272+:8] = 8'hbb;\
sBoxLayer[280+:8] = 8'hb0;\
sBoxLayer[288+:8] = 8'hb2;\
sBoxLayer[296+:8] = 8'hb1;\
sBoxLayer[304+:8] = 8'hb4;\
sBoxLayer[312+:8] = 8'hbf;\
sBoxLayer[320+:8] = 8'hb7;\
sBoxLayer[328+:8] = 8'hba;\
sBoxLayer[336+:8] = 8'hb8;\
sBoxLayer[344+:8] = 8'hb5;\
sBoxLayer[352+:8] = 8'hb9;\
sBoxLayer[360+:8] = 8'hbc;\
sBoxLayer[368+:8] = 8'hb3;\
sBoxLayer[376+:8] = 8'hb6;\
sBoxLayer[384+:8] = 8'h0e;\
sBoxLayer[392+:8] = 8'h0d;\
sBoxLayer[400+:8] = 8'h0b;\
sBoxLayer[408+:8] = 8'h00;\
sBoxLayer[416+:8] = 8'h02;\
sBoxLayer[424+:8] = 8'h01;\
sBoxLayer[432+:8] = 8'h04;\
sBoxLayer[440+:8] = 8'h0f;\
sBoxLayer[448+:8] = 8'h07;\
sBoxLayer[456+:8] = 8'h0a;\
sBoxLayer[464+:8] = 8'h08;\
sBoxLayer[472+:8] = 8'h05;\
sBoxLayer[480+:8] = 8'h09;\
sBoxLayer[488+:8] = 8'h0c;\
sBoxLayer[496+:8] = 8'h03;\
sBoxLayer[504+:8] = 8'h06;\
sBoxLayer[512+:8] = 8'h2e;\
sBoxLayer[520+:8] = 8'h2d;\
sBoxLayer[528+:8] = 8'h2b;\
sBoxLayer[536+:8] = 8'h20;\
sBoxLayer[544+:8] = 8'h22;\
sBoxLayer[552+:8] = 8'h21;\
sBoxLayer[560+:8] = 8'h24;\
sBoxLayer[568+:8] = 8'h2f;\
sBoxLayer[576+:8] = 8'h27;\
sBoxLayer[584+:8] = 8'h2a;\
sBoxLayer[592+:8] = 8'h28;\
sBoxLayer[600+:8] = 8'h25;\
sBoxLayer[608+:8] = 8'h29;\
sBoxLayer[616+:8] = 8'h2c;\
sBoxLayer[624+:8] = 8'h23;\
sBoxLayer[632+:8] = 8'h26;\
sBoxLayer[640+:8] = 8'h1e;\
sBoxLayer[648+:8] = 8'h1d;\
sBoxLayer[656+:8] = 8'h1b;\
sBoxLayer[664+:8] = 8'h10;\
sBoxLayer[672+:8] = 8'h12;\
sBoxLayer[680+:8] = 8'h11;\
sBoxLayer[688+:8] = 8'h14;\
sBoxLayer[696+:8] = 8'h1f;\
sBoxLayer[704+:8] = 8'h17;\
sBoxLayer[712+:8] = 8'h1a;\
sBoxLayer[720+:8] = 8'h18;\
sBoxLayer[728+:8] = 8'h15;\
sBoxLayer[736+:8] = 8'h19;\
sBoxLayer[744+:8] = 8'h1c;\
sBoxLayer[752+:8] = 8'h13;\
sBoxLayer[760+:8] = 8'h16;\
sBoxLayer[768+:8] = 8'h4e;\
sBoxLayer[776+:8] = 8'h4d;\
sBoxLayer[784+:8] = 8'h4b;\
sBoxLayer[792+:8] = 8'h40;\
sBoxLayer[800+:8] = 8'h42;\
sBoxLayer[808+:8] = 8'h41;\
sBoxLayer[816+:8] = 8'h44;\
sBoxLayer[824+:8] = 8'h4f;\
sBoxLayer[832+:8] = 8'h47;\
sBoxLayer[840+:8] = 8'h4a;\
sBoxLayer[848+:8] = 8'h48;\
sBoxLayer[856+:8] = 8'h45;\
sBoxLayer[864+:8] = 8'h49;\
sBoxLayer[872+:8] = 8'h4c;\
sBoxLayer[880+:8] = 8'h43;\
sBoxLayer[888+:8] = 8'h46;\
sBoxLayer[896+:8] = 8'hfe;\
sBoxLayer[904+:8] = 8'hfd;\
sBoxLayer[912+:8] = 8'hfb;\
sBoxLayer[920+:8] = 8'hf0;\
sBoxLayer[928+:8] = 8'hf2;\
sBoxLayer[936+:8] = 8'hf1;\
sBoxLayer[944+:8] = 8'hf4;\
sBoxLayer[952+:8] = 8'hff;\
sBoxLayer[960+:8] = 8'hf7;\
sBoxLayer[968+:8] = 8'hfa;\
sBoxLayer[976+:8] = 8'hf8;\
sBoxLayer[984+:8] = 8'hf5;\
sBoxLayer[992+:8] = 8'hf9;\
sBoxLayer[1000+:8] = 8'hfc;\
sBoxLayer[1008+:8] = 8'hf3;\
sBoxLayer[1016+:8] = 8'hf6;\
sBoxLayer[1024+:8] = 8'h7e;\
sBoxLayer[1032+:8] = 8'h7d;\
sBoxLayer[1040+:8] = 8'h7b;\
sBoxLayer[1048+:8] = 8'h70;\
sBoxLayer[1056+:8] = 8'h72;\
sBoxLayer[1064+:8] = 8'h71;\
sBoxLayer[1072+:8] = 8'h74;\
sBoxLayer[1080+:8] = 8'h7f;\
sBoxLayer[1088+:8] = 8'h77;\
sBoxLayer[1096+:8] = 8'h7a;\
sBoxLayer[1104+:8] = 8'h78;\
sBoxLayer[1112+:8] = 8'h75;\
sBoxLayer[1120+:8] = 8'h79;\
sBoxLayer[1128+:8] = 8'h7c;\
sBoxLayer[1136+:8] = 8'h73;\
sBoxLayer[1144+:8] = 8'h76;\
sBoxLayer[1152+:8] = 8'hae;\
sBoxLayer[1160+:8] = 8'had;\
sBoxLayer[1168+:8] = 8'hab;\
sBoxLayer[1176+:8] = 8'ha0;\
sBoxLayer[1184+:8] = 8'ha2;\
sBoxLayer[1192+:8] = 8'ha1;\
sBoxLayer[1200+:8] = 8'ha4;\
sBoxLayer[1208+:8] = 8'haf;\
sBoxLayer[1216+:8] = 8'ha7;\
sBoxLayer[1224+:8] = 8'haa;\
sBoxLayer[1232+:8] = 8'ha8;\
sBoxLayer[1240+:8] = 8'ha5;\
sBoxLayer[1248+:8] = 8'ha9;\
sBoxLayer[1256+:8] = 8'hac;\
sBoxLayer[1264+:8] = 8'ha3;\
sBoxLayer[1272+:8] = 8'ha6;\
sBoxLayer[1280+:8] = 8'h8e;\
sBoxLayer[1288+:8] = 8'h8d;\
sBoxLayer[1296+:8] = 8'h8b;\
sBoxLayer[1304+:8] = 8'h80;\
sBoxLayer[1312+:8] = 8'h82;\
sBoxLayer[1320+:8] = 8'h81;\
sBoxLayer[1328+:8] = 8'h84;\
sBoxLayer[1336+:8] = 8'h8f;\
sBoxLayer[1344+:8] = 8'h87;\
sBoxLayer[1352+:8] = 8'h8a;\
sBoxLayer[1360+:8] = 8'h88;\
sBoxLayer[1368+:8] = 8'h85;\
sBoxLayer[1376+:8] = 8'h89;\
sBoxLayer[1384+:8] = 8'h8c;\
sBoxLayer[1392+:8] = 8'h83;\
sBoxLayer[1400+:8] = 8'h86;\
sBoxLayer[1408+:8] = 8'h5e;\
sBoxLayer[1416+:8] = 8'h5d;\
sBoxLayer[1424+:8] = 8'h5b;\
sBoxLayer[1432+:8] = 8'h50;\
sBoxLayer[1440+:8] = 8'h52;\
sBoxLayer[1448+:8] = 8'h51;\
sBoxLayer[1456+:8] = 8'h54;\
sBoxLayer[1464+:8] = 8'h5f;\
sBoxLayer[1472+:8] = 8'h57;\
sBoxLayer[1480+:8] = 8'h5a;\
sBoxLayer[1488+:8] = 8'h58;\
sBoxLayer[1496+:8] = 8'h55;\
sBoxLayer[1504+:8] = 8'h59;\
sBoxLayer[1512+:8] = 8'h5c;\
sBoxLayer[1520+:8] = 8'h53;\
sBoxLayer[1528+:8] = 8'h56;\
sBoxLayer[1536+:8] = 8'h9e;\
sBoxLayer[1544+:8] = 8'h9d;\
sBoxLayer[1552+:8] = 8'h9b;\
sBoxLayer[1560+:8] = 8'h90;\
sBoxLayer[1568+:8] = 8'h92;\
sBoxLayer[1576+:8] = 8'h91;\
sBoxLayer[1584+:8] = 8'h94;\
sBoxLayer[1592+:8] = 8'h9f;\
sBoxLayer[1600+:8] = 8'h97;\
sBoxLayer[1608+:8] = 8'h9a;\
sBoxLayer[1616+:8] = 8'h98;\
sBoxLayer[1624+:8] = 8'h95;\
sBoxLayer[1632+:8] = 8'h99;\
sBoxLayer[1640+:8] = 8'h9c;\
sBoxLayer[1648+:8] = 8'h93;\
sBoxLayer[1656+:8] = 8'h96;\
sBoxLayer[1664+:8] = 8'hce;\
sBoxLayer[1672+:8] = 8'hcd;\
sBoxLayer[1680+:8] = 8'hcb;\
sBoxLayer[1688+:8] = 8'hc0;\
sBoxLayer[1696+:8] = 8'hc2;\
sBoxLayer[1704+:8] = 8'hc1;\
sBoxLayer[1712+:8] = 8'hc4;\
sBoxLayer[1720+:8] = 8'hcf;\
sBoxLayer[1728+:8] = 8'hc7;\
sBoxLayer[1736+:8] = 8'hca;\
sBoxLayer[1744+:8] = 8'hc8;\
sBoxLayer[1752+:8] = 8'hc5;\
sBoxLayer[1760+:8] = 8'hc9;\
sBoxLayer[1768+:8] = 8'hcc;\
sBoxLayer[1776+:8] = 8'hc3;\
sBoxLayer[1784+:8] = 8'hc6;\
sBoxLayer[1792+:8] = 8'h3e;\
sBoxLayer[1800+:8] = 8'h3d;\
sBoxLayer[1808+:8] = 8'h3b;\
sBoxLayer[1816+:8] = 8'h30;\
sBoxLayer[1824+:8] = 8'h32;\
sBoxLayer[1832+:8] = 8'h31;\
sBoxLayer[1840+:8] = 8'h34;\
sBoxLayer[1848+:8] = 8'h3f;\
sBoxLayer[1856+:8] = 8'h37;\
sBoxLayer[1864+:8] = 8'h3a;\
sBoxLayer[1872+:8] = 8'h38;\
sBoxLayer[1880+:8] = 8'h35;\
sBoxLayer[1888+:8] = 8'h39;\
sBoxLayer[1896+:8] = 8'h3c;\
sBoxLayer[1904+:8] = 8'h33;\
sBoxLayer[1912+:8] = 8'h36;\
sBoxLayer[1920+:8] = 8'h6e;\
sBoxLayer[1928+:8] = 8'h6d;\
sBoxLayer[1936+:8] = 8'h6b;\
sBoxLayer[1944+:8] = 8'h60;\
sBoxLayer[1952+:8] = 8'h62;\
sBoxLayer[1960+:8] = 8'h61;\
sBoxLayer[1968+:8] = 8'h64;\
sBoxLayer[1976+:8] = 8'h6f;\
sBoxLayer[1984+:8] = 8'h67;\
sBoxLayer[1992+:8] = 8'h6a;\
sBoxLayer[2000+:8] = 8'h68;\
sBoxLayer[2008+:8] = 8'h65;\
sBoxLayer[2016+:8] = 8'h69;\
sBoxLayer[2024+:8] = 8'h6c;\
sBoxLayer[2032+:8] = 8'h63;\
sBoxLayer[2040+:8] = 8'h66;
`endif